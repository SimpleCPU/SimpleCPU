// Exception Unit
module exception_unit ();

endmodule
