library verilog;
use verilog.vl_types.all;
entity top_tb is
end top_tb;
