module exception_unit ();

endmodule
