// Exception Unit
// Work in progress
module exception_unit ();

endmodule
