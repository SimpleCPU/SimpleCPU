library verilog;
use verilog.vl_types.all;
entity boot_code_sv_unit is
end boot_code_sv_unit;
