library verilog;
use verilog.vl_types.all;
entity init_imem_sv_unit is
end init_imem_sv_unit;
