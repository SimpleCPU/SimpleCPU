// Memory initialisation

function void init_imem ();
    T1.I_MEM1.imem [0] = 32'h10000011;
    T1.I_MEM1.imem [1] = 32'h10000011;
    T1.I_MEM1.imem [2] = 32'h20000022;
    T1.I_MEM1.imem [3] = 32'h30000033;
    T1.I_MEM1.imem [4] = 32'h40000044;
    T1.I_MEM1.imem [5] = 32'h50000055;
    T1.I_MEM1.imem [6] = 32'h60000066;
    T1.I_MEM1.imem [7] = 32'h70000077;
    T1.I_MEM1.imem [8] = 32'h80000088;
    T1.I_MEM1.imem [9] = 32'h90000099;

endfunction
