// Top module connecting all the other modules

module top
    (
        input   wire    clk,
        input   wire    reset
    );

endmodule
