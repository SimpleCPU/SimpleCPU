library verilog;
use verilog.vl_types.all;
entity init_dmem_sv_unit is
end init_dmem_sv_unit;
